* AD8512 SPICE Macro-model                   
* Description: Amplifier
* Generic Desc: 10/30V, JFET, OP, Low Noise, Low Ib, 2X
* Developed by: GEC/ADSJ
* Revision History: 08/10/2012 - Updated to new header style
* 1.1 (08/2009)
* Copyright 2002, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes: Derived from AD8510 Rev. 1.0 SB, ADSiV apps, 04/2002
*		VSY=5V, T=25�C
*
* Not Modeled:
*    
* Parameters modeled include: 
* This model simulates typical values for the B grade AD8510
*
* END Notes
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD8512   1 2 99 50 30
*
* INPUT STAGE
*
R3   5  50    3.385E3
R4   6  50   3.385E3
CIN  1   2    5.5E-12
I1     99  4  2.954E-4
V10   4     55 DC 4
D10  55   99 DX
IOS  1   2    6E-12
EOS  60  1    POLY(2)  (17, 24) (73, 24)  80E-6  1 1
EN   7  60    42  0  1
GN1  0   1    45  0  1E-6
GN2  0   2    48  0  1E-6
J1   5   2    4   JX
J2   6   7    4   JX
GB1  2  50    POLY(3) (4, 2) (5, 2) (50, 2) 1E-12 1E-12 1E-12
GB2  7  50    POLY(3) (4, 7) (6, 7) (50, 7) 1E-12 1E-12 1E-12
*
EREF 98  0    24  0   1
*
* VOLTAGE NOISE GENERATOR
*
VN1  41  0    DC 2
DN1  41 42    DEN
DN2  42 43    DEN
VN2  0  43    DC 2
*
* CURRENT NOISE GENERATOR
*
VN3  44  0    DC 2
DN3  44 45    DIN
DN4  45 46    DIN
VN4  0  46    DC 2
*
* CURRENT NOISE GENERATOR
*
VN5  47  0    DC 2
DN5  47 48    DIN
DN6  48 49    DIN
VN6  0  49    DC 2
*  
* SECOND STAGE & POLE AT 50 Hz
*
R5   9  98  8.16E4
C3   9  98    39E-9
G1   98  9    5  6  7.8E-1
V2   99  8    1.8
V3   10 50   1.8
D1   9   8    DX
D2   10  9    DX
*
* CMRR WITH ZERO AT 297 Hz
*
R11  16 17     8E+06
C8   16 17     6.695E-11
R12  17  98    8
E3   16 98     POLY(2) (98, 2)  (98, 0)  1.00 1.00
*
* PSRR WITH ZERO AT 0.5 Hz
*
EPSY 72 98 POLY(1) (99,50) 0 5
CPS3 72 73 1E-9
RPS3 72 73 316.2E+6
RPS4 73 98 1
*
* POLE AT 13.8 MHZ
*
R13  18 98     1E3
C9   18 98    11.5E-12
G5   98 18     9  24  1E-3
*
* OUTPUT STAGE
*
R14  24 99     500E3
R15  24 50     500E3
CF   24  0     1E-6
ISY  99 50     1.9E-3
R16  29 99     180
R17  29 50     180
L1    29 30     1E-8
G6   27 50     18 29  9.09E-3
G7   28 50     29 18  9.09E-3
G8   29 99     99 18  5.5555E-03
G9   50 29     18 50  5.5555E-03
V4   25 29     6.675
V5   29 26     6.675
D3   18 25     DX
D4   26 18     DX
D5   99 27     DX
D6   99 28     DX
D7   50 27     DY
D8   50 28     DY
F1   29  0     V4  1
F2   0  29     V5  1
*
* MODELS USED
*
.MODEL JX PJF(BETA=1.4E-3 VTO=-1.00  IS=75E-12 RD=0
+ RS=0 CGD=1E-12 CGS=1E-12)
.MODEL DX   D(IS=1E-15 RS=0 CJO=1E-12)
.MODEL DY   D(IS=1E-15 BV=50 RS=10 CJO=1E-12)
.MODEL DEN  D(IS=1E-12, RS=3400, KF=0.35E-14, AF=0.830)
.MODEL DIN  D(IS=1E-12, RS=19.3E-6, KF=4.28E-15, AF=1)
.ENDS AD8512






