PIEZO AMP

.inc third-party/ad8512.cir
.inc third-party/lm358.lib

* power
VCC hardvcc gnd DC 10
R1 hardvcc vcc 1

* voltage divider
R2 vcc halfu 10k
R3 halfu gnd 10k

* middle voltage buffer
xop1 halfu half vcc gnd half ad8512
chalf half gnd 10u

*generator
*vin signal gnd DC 5.25

* generator
*Csingnal signal1 signal 20n
*Rsignal signal0 signal1 1
VGEN signal0 half SIN(1 0.1 50)
*VGEN signal0 half PWL(0ms 0 1ms 1 2ms 0 3ms -1 4ms 0 5ms 0) r=0
*VGEN signal0 half PWL(0ms 0 10ms 0.05 20ms 0 40ms 0) r=0
*VGEN signal0 half PWL(0ms 0 1ms 0 1ms 1 2ms 1 2ms 0 4ms 0) r=0
VGEN signal0 half PWL(0s 0 0.2s 0 0.2s 0.2 0.4s 0.2 0.4s 0 0.6s 0) r=0

xamp signal vcc half gnd out ina amplifier

.subckt amplifier input vcc mid gnd output input_amp
rz1 input gnd 1000K
rz2 input vcc 1000K
xpreamp input input_amp vcc gnd input_amp lm358
*cpreamp input_amp0 input_amp 10u
xop mid in- vcc gnd output lm358
*r3 input_amp gnd 200K
*r4 input_amp vcc 200K
r0 input_amp in- 7K
c in- output 6u
r in- output 250K
.ends

.control
    tran 0.01ms 1500ms 100ms
    plot V(signal) V(out) 
.endc
.end
