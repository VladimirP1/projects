PIEZO AMP

.inc third-party/ad8512.cir
.inc third-party/lm358.lib

* power
VCC hardvcc gnd DC 10
R1 hardvcc vcc 1

* voltage divider
R2 vcc halfu 10k
R3 halfu gnd 10k

* middle voltage buffer
xop1 halfu half vcc gnd half ad8512
chalf half gnd 10u

* generator
Csingnal signal1 signal 200u
Rsignal signal0 signal1 1
*VGEN signal0 half SIN(1 0.1 50)
*VGEN signal0 half PWL(0ms 0 1ms 1 2ms 0 3ms -1 4ms 0 5ms 0) r=0
*VGEN signal0 half PWL(0ms 0 10ms 0.05 20ms 0 40ms 0) r=0
*VGEN signal0 half PWL(0ms 0 1ms 0 1ms 1 2ms 1 2ms 0 4ms 0) r=0
VGEN signal0 half PWL(0s 0 0.2s 0 0.2s 0.2 0.4s 0.2 0.4s 0 1s 0) r=0

xamp signal vcc half gnd out ina amplifier

.subckt amplifier input vcc mid gnd output input_amp 
cpreamp input input_amp 100u ic=0v
xop mid in- vcc gnd output ad8512
r0 input_amp in- 7K
c1 in- output 6u
r1 in- output 250K
*r2 input_amp output 10meg
.ends

.control
    tran 2ms 10000ms 500ms uic
    plot V(signal) V(out) V(ina)
.endc
.end
