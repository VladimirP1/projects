VOLTAGE DIVIDER

.inc third-party/lm358.lib
.inc third-party/ad8512.cir
* power
VCC hardvcc gnd DC 10
R1 hardvcc vcc 1

* voltage divider
R2 vcc halfu 10k
R3 halfu gnd 10k

* middle voltage buffer
xop1 halfu half vcc gnd half ad8512
chalf half gnd 10u

* generator
VGEN signal half SIN(0 0.1 10K)


xamp signal vcc half gnd out amplifier

.subckt amplifier input vcc mid gnd output
xopa mid inrc vcc gnd output ad8512
R0 input inputr 0
C1 inputr inrc 0.01u
R1 inrc output 1K
*C2 inrc output 0.001u
.ends

.control
    tran 10ns 1ms
    plot V(signal) V(out) V(half)
.endc
.end
